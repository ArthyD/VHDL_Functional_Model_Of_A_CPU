library work;
use work.bit_vector_natural_pack.all;


entity Test is
end Test;

architecture bit_vector_natural_pack_test of Test is
begin
    process
        constant test_bit_vector: bit_vector <= "11001100"; -- 0b11001100 is dec(204)
        constant test_data_width: natural <= 8; -- 0b11001100 are 8 bits
        constant test_integer: integer <= 204; -- dec(204) is 0b11001100
        
        constant converted_integer <= bit_vector2natural(test_bit_vector);
        constant converted_bit_vector <= natural2bit_vector(test_integer, test_data_width);

        assert test_bit_vector == converted_bit_vector;
        assert test_integer == converted_integer;
    end process
end architecture
